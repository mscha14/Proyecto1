`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// Estudents: Mauricio Salomón----Michael Chaves
// 
// Create Date:    16:41:29 07/30/2015 
// Design Name: 
// Module Name:   MEM_uPROGRAMA
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: //memoria microprogramada, contiene todas las instrucciones de la máquina de estados.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module MEM_uPROGRAMA(DIR, SALIDAS);

	input [4:0] DIR;
	output reg [21:0] SALIDAS;

	always @ (DIR)
	case(DIR)

			5'b00000:	SALIDAS = 22'b001_00000_1001111_1110_000;
			5'b00001:	SALIDAS = 22'b010_00111_0010010_1110_000;
			5'b00010:	SALIDAS = 22'b011_10110_0000110_1110_000;
			5'b00011:	SALIDAS = 22'b100_11101_1001100_1110_000;
			5'b00100:	SALIDAS = 22'b001_00000_0100100_1110_000;
			5'b00101:	SALIDAS = 22'b101_00001_0100100_1110_000;
			5'b00110:	SALIDAS = 22'b000_00101_0100100_1110_000;
			5'b00111:	SALIDAS = 22'b001_00000_0010010_1110_011;
			5'b01000:	SALIDAS = 22'b011_01100_0100000_1110_011;
			5'b01001:	SALIDAS = 22'b100_10011_0001111_1110_011;
			5'b01010:	SALIDAS = 22'b101_00001_0100100_1110_011;
			5'b01011:	SALIDAS = 22'b000_01010_0100100_1110_011;
			5'b01100:	SALIDAS = 22'b001_00000_0100000_1110_101;
			5'b01101:	SALIDAS = 22'b100_10000_0000000_1110_101;
			5'b01110:	SALIDAS = 22'b101_00001_0100100_1110_101;
			5'b01111:	SALIDAS = 22'b000_01110_0100100_1110_101;
			5'b10000:	SALIDAS = 22'b001_00000_0000000_1110_001;
			5'b10001:	SALIDAS = 22'b101_00001_0100100_1110_001;
			5'b10010:	SALIDAS = 22'b000_10001_0100100_1110_001;
			5'b10011:	SALIDAS = 22'b001_00000_0001111_1110_001;
			5'b10100:	SALIDAS = 22'b101_00001_0100100_1110_001;
			5'b10101:	SALIDAS = 22'b000_10100_0100100_1110_001;
			5'b10110:	SALIDAS = 22'b001_00000_0000110_1110_001;
			5'b10111:	SALIDAS = 22'b100_11010_0001100_1110_001;
			5'b11000:	SALIDAS = 22'b101_00001_0100100_1110_001;
			5'b11001:	SALIDAS = 22'b000_11000_0100100_1110_001;
			5'b11010:	SALIDAS = 22'b001_00000_0001100_1110_001;
			5'b11011:	SALIDAS = 22'b101_00001_0100100_1110_001;
			5'b11100:	SALIDAS = 22'b000_11011_0100100_1110_001;
			5'b11101:	SALIDAS = 22'b001_00000_1001100_1110_001;
			5'b11110:	SALIDAS = 22'b000_11011_1001100_1110_001;
			
			
		default:	SALIDAS = 22'b001_00000_1001111_1110_000;

		endcase


endmodule
